
library ieee;
use ieee.std_logic_1164.all;

entity tb_float is
  port (
    ok   : out std_ulogic;
    done : out std_ulogic);
end entity tb_float;

library work;
use work.float.float32;

architecture behavior of tb_float is

begin

  

end architecture behavior;
